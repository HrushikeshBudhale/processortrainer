//Width related constant
`define INAT_WIDTH 32
`define REG_ADDR_WIDTH 5
`define LITERAL_WIDTH 16
//Opcode 
`define ADD 8'h20
`define ADDC 8'h30
`define AND 8'h28
`define ANDC 8'h38
`define BEQ 8h'1D
`define BNE 8'h1E
`define COMPEQ 8'h24
`define COMPEQC 8'h34
`define CMPLE 8'h26
`define CMPLEC 8'h36
`define CMPLT 8'h25
`define CMPLTC 8'h35
`define DIV 8'h23
`define DIVC 8'h33
`define JMP 8'h1B
`define L 8'h18
`define LDR 8'h1F
`define MUL	8'h22
`define MULC 8'h32
`define OR 8'h29
`define ORC 8'h39
`define SHL	8'h2C
`define SHLC 8'h3C
`define SHR 8'h2D
`define SHRC 8'h3D
`define SRA 8'h2E
`define SRAC 8'h3E
`define SUB 8'h21
`define SUBC 8'h21
`define ST 8'h19
`define XOR 8'h2A
`define XORC 8'h3A
//ALU OPCODE 
`define ALU_ADD 8'h00
`define ALU_SUB 8'h01
`define ALU_AND 8'h18
`define ALU_OR 8'h1E
`define ALU_XOR 8'h16
`define ALU_LDR 8'h1A
`define ALU_SHL 8'h20
`define ALU_SHR 8'h21
`define ALU_SRA 8'h23
`define ALU_CMPEQ 8'h33
`define ALU_CMPLT 8'h35
`define ALU_CMPLE 8'h37
`define ALU_MUL 8'h02
`define ALU_DIV 8'h03
